`timescale 10 ns / 1 ns

module mul(
	input clk,
	input rst,
	input [31:0] a,
	input [31:0] b,
	input valid,
	output ready,
	output [63:0] result
);

endmodule
